method module_l3_switch_forward_table_add_entry=ingress.module_l3_switch_forward_table_add_entry;
method module_l3_switch_ipv4_nhop_add_entry=ingress.module_l3_switch_ipv4_nhop_add_entry;
method module_l3_switch_send_frame_add_entry=ingress.module_l3_switch_send_frame_add_entry;
