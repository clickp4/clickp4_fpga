method Action module_if_if_equal_add_entry(ModuleIfIfEqualReqT key, ModuleIfIfEqualRspT val);
method Action module_if_if_large_add_entry(ModuleIfIfLargeReqT key, ModuleIfIfLargeRspT val);
method Action module_if_if_small_add_entry(ModuleIfIfSmallReqT key, ModuleIfIfSmallRspT val);
method Action pipeline_start_tbl_pipeline_start_add_entry(PipelineStartTblPipelineStartReqT key, PipelineStartTblPipelineStartRspT val);
