import Ethernet::*;
import StructDefines::*;
typedef union tagged {
    struct {
    } ReqT;
    struct {
    } ReqT;
} ModuleIfIfEqualParam deriving (Bits, Eq, FShow);
typedef union tagged {
    struct {
    } ReqT;
    struct {
    } ReqT;
} ModuleIfIfLargeParam deriving (Bits, Eq, FShow);
typedef union tagged {
    struct {
    } ReqT;
    struct {
    } ReqT;
} ModuleIfIfSmallParam deriving (Bits, Eq, FShow);
import Ethernet::*;
import StructDefines::*;
