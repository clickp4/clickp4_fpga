method module_if_if_equal_add_entry = prog.module_if_if_equal_add_entry;
method module_if_if_large_add_entry = prog.module_if_if_large_add_entry;
method module_if_if_small_add_entry = prog.module_if_if_small_add_entry;
method pipeline_start_tbl_pipeline_start_add_entry = prog.pipeline_start_tbl_pipeline_start_add_entry;
