import Ethernet::*;
import StructDefines::*;
typedef union tagged {
    struct {
    } ReqT;
    struct {
    } ReqT;
} ModuleForForEndParam deriving (Bits, Eq, FShow);
typedef union tagged {
    struct {
    } ReqT;
    struct {
    } ReqT;
} ModuleForForInitParam deriving (Bits, Eq, FShow);
typedef union tagged {
    struct {
    } ReqT;
    struct {
    } ReqT;
} ModuleForForLoopParam deriving (Bits, Eq, FShow);
import Ethernet::*;
import StructDefines::*;
