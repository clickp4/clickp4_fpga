method Action pipeline_rewind_rewind_table_add_entry(PipelineRewindRewindTableReqT key, PipelineRewindRewindTableRspT val);
