method module_if_if_equal_add_entry = prog.module_if_if_equal_add_entry;
method module_if_if_large_add_entry = prog.module_if_if_large_add_entry;
method module_if_if_small_add_entry = prog.module_if_if_small_add_entry;
