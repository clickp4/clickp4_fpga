method pipeline_start_tbl_pipeline_start_add_entry=ingress.pipeline_start_tbl_pipeline_start_add_entry;
