import Ethernet::*;
import StructDefines::*;
typedef union tagged {
    struct {
    } ReqT;
    struct {
    } ReqT;
} PipelineRewindRewindTableParam deriving (Bits, Eq, FShow);
import Ethernet::*;
import StructDefines::*;
