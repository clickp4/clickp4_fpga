`define PARSER Parser
`define DEPARSER Deparser
`define MATCHTABLE Control
`define TYPEDEF StructDefines
`define NUM_RXCHAN 1
`define NUM_TXCHAN 1
`define NUM_HOSTCHAN 1
`define STREAM 
`define NUM_RXCHAN 1
`define NUM_TXCHAN 1
`define NUM_HOSTCHAN 1
`define NUM_METAGEN 1
`define NUM_PKTGEN 1
`define STREAM 
`define NicVersion 1579743661
`define DataBusWidth 128
`define IMPORT_HOSTIF 
`define BYTE_ENABLES 
`define ClockDefaultParam 
`define ConnectalVersion 16.11.1
`define NumberOfMasters 1
`define PinType Empty
`define PinTypeInclude Misc
`define NumberOfUserTiles 1
`define SlaveDataBusWidth 32
`define SlaveControlAddrWidth 5
`define BurstLenSize 12
`define project_dir $(DTOP)
`define MainClockPeriod 20
`define DerivedClockPeriod 10.000000
`define CnocTop 
`define XsimHostInterface 
`define PhysAddrWidth 40
`define SIMULATION 
`define CONNECTAL_BITS_DEPENDENCES bsim
`define BOARD_bluesim 
