method Action module_firewall_firewall_with_tcp_add_entry(ModuleFirewallFirewallWithTcpReqT key, ModuleFirewallFirewallWithTcpRspT val);
method Action module_firewall_firewall_with_udp_add_entry(ModuleFirewallFirewallWithUdpReqT key, ModuleFirewallFirewallWithUdpRspT val);
