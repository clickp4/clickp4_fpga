method module_if_if_equal_add_entry=ingress.module_if_if_equal_add_entry;
method module_if_if_large_add_entry=ingress.module_if_if_large_add_entry;
method module_if_if_small_add_entry=ingress.module_if_if_small_add_entry;
