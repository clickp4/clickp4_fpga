method module_firewall_firewall_with_tcp_add_entry=ingress.module_firewall_firewall_with_tcp_add_entry;
method module_firewall_firewall_with_udp_add_entry=ingress.module_firewall_firewall_with_udp_add_entry;
method pipeline_start_tbl_pipeline_start_add_entry=ingress.pipeline_start_tbl_pipeline_start_add_entry;
