import Ethernet::*;
import StructDefines::*;
typedef union tagged {
    struct {
    } ReqT;
    struct {
    } ReqT;
    struct {
    } ReqT;
} PipelineStartTblPipelineStartParam deriving (Bits, Eq, FShow);
import Ethernet::*;
import StructDefines::*;
