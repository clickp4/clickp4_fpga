`define PARSER Parser
`define DEPARSER Deparser
`define MATCHTABLE Control
`define TYPEDEF StructDefines
`define NUM_RXCHAN 1
`define NUM_TXCHAN 1
`define NUM_HOSTCHAN 1
`define STREAM 
`define NUM_RXCHAN 1
`define NUM_TXCHAN 1
`define NUM_HOSTCHAN 1
`define NUM_METAGEN 1
`define NUM_PKTGEN 1
`define STREAM 
`define NicVersion 2597774736
`define DataBusWidth 128
`define IMPORT_HOSTIF 
`define BYTE_ENABLES 
`define ClockDefaultParam 
`define XILINX_SYS_CLK 
`define ConnectalVersion 16.11.1
`define NumberOfMasters 1
`define PinType NfsumePins
`define PinTypeInclude NfsumePins
`define NumberOfUserTiles 1
`define SlaveDataBusWidth 32
`define SlaveControlAddrWidth 5
`define BurstLenSize 12
`define project_dir $(DTOP)
`define MainClockPeriod 4
`define DerivedClockPeriod 4.000000
`define PcieClockPeriod 4
`define XILINX 1
`define Virtex7 
`define PCIE 
`define PCIE3 
`define PcieHostInterface 
`define PhysAddrWidth 40
`define NUMBER_OF_LEDS 2
`define PcieLanes 8
`define CONNECTAL_BITS_DEPENDENCES hw/mkTop.bit
`define CONNECTAL_RUN_SCRIPT $(CONNECTALDIR)/scripts/run.pcietest
`define BOARD_nfsume 
