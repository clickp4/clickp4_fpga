method Action module_for_for_end_add_entry(ModuleForForEndReqT key, ModuleForForEndRspT val);
method Action module_for_for_init_add_entry(ModuleForForInitReqT key, ModuleForForInitRspT val);
method Action module_for_for_loop_add_entry(ModuleForForLoopReqT key, ModuleForForLoopRspT val);
method Action pipeline_start_tbl_pipeline_start_add_entry(PipelineStartTblPipelineStartReqT key, PipelineStartTblPipelineStartRspT val);
