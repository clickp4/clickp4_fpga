import Ethernet::*;
import StructDefines::*;
typedef union tagged {
    struct {
    } ReqT;
    struct {
    } ReqT;
    struct {
    } ReqT;
} ModuleFirewallFirewallWithTcpParam deriving (Bits, Eq, FShow);
typedef union tagged {
    struct {
    } ReqT;
    struct {
    } ReqT;
    struct {
    } ReqT;
} ModuleFirewallFirewallWithUdpParam deriving (Bits, Eq, FShow);
import Ethernet::*;
import StructDefines::*;
