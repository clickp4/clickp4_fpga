import Ethernet::*;
import StructDefines::*;
typedef union tagged {
    struct {
    } ReqT;
    struct {
    } ReqT;
} ModuleL3SwitchForwardTableParam deriving (Bits, Eq, FShow);
typedef union tagged {
    struct {
    } ReqT;
    struct {
    } ReqT;
    struct {
    } ReqT;
} ModuleL3SwitchIpv4NhopParam deriving (Bits, Eq, FShow);
typedef union tagged {
    struct {
    } ReqT;
    struct {
    } ReqT;
    struct {
    } ReqT;
} ModuleL3SwitchSendFrameParam deriving (Bits, Eq, FShow);
typedef union tagged {
    struct {
    } ReqT;
    struct {
    } ReqT;
    struct {
    } ReqT;
} PipelineStartTblPipelineStartParam deriving (Bits, Eq, FShow);
import Ethernet::*;
import StructDefines::*;
