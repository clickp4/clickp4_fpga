method module_while_while_equal_add_entry = prog.module_while_while_equal_add_entry;
method module_while_while_init_add_entry = prog.module_while_while_init_add_entry;
method module_while_while_large_add_entry = prog.module_while_while_large_add_entry;
method module_while_while_small_add_entry = prog.module_while_while_small_add_entry;
method pipeline_start_tbl_pipeline_start_add_entry = prog.pipeline_start_tbl_pipeline_start_add_entry;
