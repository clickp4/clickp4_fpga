method pipeline_rewind_rewind_table_add_entry=ingress.pipeline_rewind_rewind_table_add_entry;
