`define PARSER Parser
`define DEPARSER Deparser
`define MATCHTABLE Control
`define TYPEDEF StructDefines
`define NUM_RXCHAN 1
`define NUM_TXCHAN 1
`define NUM_HOSTCHAN 1
`define STREAM 
`define NUM_RXCHAN 1
`define NUM_TXCHAN 1
`define NUM_HOSTCHAN 1
`define NUM_METAGEN 1
`define NUM_PKTGEN 1
`define STREAM 
`define NicVersion 2597774736
`define DataBusWidth 128
`define IMPORT_HOSTIF 
`define BYTE_ENABLES 
`define ClockDefaultParam 
`define ConnectalVersion 16.11.1
`define NumberOfMasters 1
`define PinType Empty
`define PinTypeInclude Misc
`define NumberOfUserTiles 1
`define SlaveDataBusWidth 32
`define SlaveControlAddrWidth 5
`define BurstLenSize 12
`define project_dir $(DTOP)
`define MainClockPeriod 8
`define DerivedClockPeriod 4.000000
`define PcieClockPeriod 8
`define XILINX 1
`define Kintex7 
`define PCIE 
`define PCIE1 
`define PcieHostInterface 
`define PhysAddrWidth 40
`define PcieLanes 8
`define CONNECTAL_BITS_DEPENDENCES hw/mkTop.bit
`define CONNECTAL_RUN_SCRIPT $(CONNECTALDIR)/scripts/run.pcietest
`define BOARD_kc705 
